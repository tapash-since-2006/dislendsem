module twotooneMUX(y,i,s0);
    input [1:0]i;
    input s0;
    output y;

    assign y=(s0?i[1]:i[0]);
endmodule

